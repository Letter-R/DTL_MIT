
import FixedPoint::*;
import Vector::*;

Vector#(9, FixedPoint#(16,16)) c =
    cons(fromReal(-0.0124), 
    cons(fromReal(0.0),
    cons(fromReal(-0.0133),
    cons(fromReal(0.0),
    cons(fromReal(0.8181),
    cons(fromReal(0.0),
    cons(fromReal(-0.0133),
    cons(fromReal(0.0),
    cons(fromReal(-0.0124),
nil)))))))));
